library IEEE;
use IEEE.std_logic_1164.all;

entity decoder8 is
        port (
                sel : in  std_logic_vector(2 downto 0);
                o  : out std_logic_vector(7 downto 0)
        );
end decoder8;

architecture decoder8_dataflow of decoder8 is
begin

	with sel select o <=
	"00000001" when "000",
	"00000010" when "001",
	"00000100" when "010",
	"00001000" when "011",
	"00010000" when "100",
	"00100000" when "101",
	"01000000" when "110",
	"10000000" when "111",
	"XXXXXXXX" when others;
end decoder8_dataflow;
